`define GET_WIDTH(N)            \
    N < 2           ?   1   :   \
    N < 4           ?   2   :   \
    N < 8           ?   3   :   \
    N < 16          ?   4   :   \
    N < 32          ?   5   :   \
    N < 64          ?   6   :   \
    N < 128         ?   7   :   \
    N < 256         ?   8   :   \
    N < 512         ?   9   :   \
    N < 1024        ?   10  :   \
    N < 2048        ?   11  :   \
    N < 4096        ?   12  :   \
    N < 8192        ?   13  :   \
    N < 16384       ?   14  :   \
    N < 32768       ?   15  :   \
    N < 65536       ?   16  :   \
    N < 131072      ?   17  :   \
    N < 262144      ?   18  :   \
    N < 524288      ?   19  :   \
    N < 1048576     ?   20  :   \
    N < 2097152     ?   21  :   \
    N < 4194304     ?   22  :   \
    N < 8388608     ?   23  :   \
    N < 16777216    ?   24  :   \
    N < 33554432    ?   25  :   \
    N < 67108864    ?   26  :   \
    N < 134217728   ?   27  :   \
    N < 268435456   ?   28  :   \
    N < 536870912   ?   29  :   \
    N < 1073741824  ?   30  :   \
    N < 2147483648  ?   31  :   \
    32

