`define HW_RESET        0
`define INVALID_INST    8
