module mmu(
    );

    // TODO

    tlb tlb();
endmodule
