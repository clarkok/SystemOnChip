`define CP0_EPC         0       // Exception PC
`define CP0_ECAUSE      1       // Exception cause
`define CP0_IE          2       // Interrupt enable
`define CP0_IS          3       // Interrupt status
`define CP0_EHB         4       // Exception handler base
`define CP0_PTB         5       // Page table base
`define CP0_PFA         6       // Page fault addr
