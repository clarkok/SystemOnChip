`define HW_RESET        0
`define MMU_PAGE_FAULT  1
`define PS2_INT         2
`define VGA_INT         3
`define UART_INT        4
`define TIMER_INT       5

`define UNALIGNED_INST  8
`define UNALIGNED_DATA  9
`define UNDEFINED_INST  10
`define PRIVILEGE_INST  11
`define PRIVILEGE_ADDR  12
`define OVERFLOW        13
`define SYSCALL         14
`define BREAK           15
